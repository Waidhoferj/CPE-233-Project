module GyroFsm (
    begin_transmission,
    recieved_data,
		end_transmission,
		clk,
		rst,
		start,
		slave_select,
		send_data,
		x_axis_data,
		y_axis_data,
		z_axis_data
);
    
endmodule